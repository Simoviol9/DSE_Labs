------------------------------------
-- Group 8 - Laboratory 6
-- Simple digital filter
-- VHDL code of memory
------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity memory is
	port (
		CLK, CS, WR, RD      : in  STD_LOGIC;
		ADDRESS  : in  STD_LOGIC_VECTOR(9 downto 0);
		DATA_IN  : in  signed(7 downto 0);
		DATA_OUT : out signed(7 downto 0));
end memory;

architecture bahaviour of memory is
	-- Define a new type variable for memory
	type mem_array is array(0 to 1023) of signed(7 downto 0);
	signal mem : mem_array := (others => (others => '0'));

	signal INTEGER_ADDRESS: INTEGER;

begin
	-- Compute the integer value of address
	INTEGER_ADDRESS <= to_integer(unsigned(ADDRESS));

	process (CLK)
	begin
		-- Writing operation (synchronous)
		if rising_edge(CLK) then
			if CS = '1' and WR = '1' then
				mem(INTEGER_ADDRESS) <= DATA_IN;
			end if;
		end if;
	end process;

	-- Reading operation (asynchronous)
	DATA_OUT <= mem(INTEGER_ADDRESS) when (CS = '1' and RD = '1') else
		(others => 'Z');
end bahaviour;
