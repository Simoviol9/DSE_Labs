-- File Part2.vhd
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
ENTITY part2 IS
	PORT (
		SW : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		HEX0, HEX1, HEX2, HEX3, HEX4 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
END part2;

ARCHITECTURE Behavior OF part2 IS
	COMPONENT mux IS
		PORT (
			SEL : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			OUTPUT : OUT STD_LOGIC_VECTOR(14 DOWNTO 0)
		);
	END COMPONENT;
	COMPONENT shifter IS
		PORT (
			INPUT : IN STD_LOGIC_VECTOR(14 DOWNTO 0);
			SEL: IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			OUTPUT : OUT STD_LOGIC_VECTOR(14 DOWNTO 0)
		);
	END COMPONENT;
	COMPONENT decoder7
		PORT (
			C : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
			DISPLAY : OUT STD_LOGIC_VECTOR(0 TO 6)
		);
	END COMPONENT;
	SIGNAL A1, A2 : STD_LOGIC_VECTOR(14 DOWNTO 0);
BEGIN
	MUX0 : mux
	PORT MAP(SW(1 DOWNTO 0), A1);
	SHIFT0 : shifter
	PORT MAP(A1, SW(4 DOWNTO 2), A2);
	H0 : decoder7
	PORT MAP(A2(2 DOWNTO 0), HEX0);
	H1 : decoder7
	PORT MAP(A2(5 DOWNTO 3), HEX1);
	H2 : decoder7
	PORT MAP(A2(8 DOWNTO 6), HEX2);
	H3 : decoder7
	PORT MAP(A2(11 DOWNTO 9), HEX3);
	H4 : decoder7
	PORT MAP(A2(14 DOWNTO 12), HEX4);
END Behavior;