LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY shifter IS
	PORT (
		INPUT : IN STD_LOGIC_VECTOR(14 DOWNTO 0);
		SEL : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
		OUTPUT : OUT STD_LOGIC_VECTOR(14 DOWNTO 0)
	);
END shifter;
ARCHITECTURE Behavior OF shifter IS
BEGIN
	PROCESS (SEL, INPUT)
	BEGIN
		IF SEL = "000" THEN
			OUTPUT <= INPUT;
		ELSIF SEL = "001" THEN
			OUTPUT(14 DOWNTO 3) <= INPUT(11 DOWNTO 0);
			OUTPUT(2 DOWNTO 0) <= INPUT(14 DOWNTO 12);
		ELSIF SEL = "010" THEN
			OUTPUT(14 DOWNTO 6) <= INPUT(8 DOWNTO 0);
			OUTPUT(5 DOWNTO 0) <= INPUT(14 DOWNTO 9);
		ELSIF SEL = "011" THEN
			OUTPUT(14 DOWNTO 9) <= INPUT(5 DOWNTO 0);
			OUTPUT(8 DOWNTO 0) <= INPUT(14 DOWNTO 6);
		ELSIF SEL = "100" THEN
			OUTPUT(14 DOWNTO 12) <= INPUT(2 DOWNTO 0);
			OUTPUT(11 DOWNTO 0) <= INPUT(14 DOWNTO 3);
		ELSE
			OUTPUT <= INPUT;
		END IF;
	END PROCESS;
END Behavior;