LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

-- Testbench for the 7 segment decoder
ENTITY part2_tb IS
END part2_tb;

ARCHITECTURE Behavior OF part2_tb IS

	COMPONENT part2
		PORT (
		SW : IN STD_LOGIC_VECTOR(4 DOWNTO 0);
		HEX0, HEX1, HEX2, HEX3, HEX4 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
	);
	END COMPONENT;

	SIGNAL DIGIT_SELECTION : STD_LOGIC_VECTOR(1 DOWNTO 0);
	SIGNAL SHIFT_SELECTION : STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL DIG0,DIG1,DIG2,DIG3,DIG4 : STD_LOGIC_VECTOR(6 DOWNTO 0);

BEGIN
	PROCESS
	BEGIN

		DIGIT_SELECTION <= "00";
		SHIFT_SELECTION <= "000";
		WAIT FOR 20 ns;
		DIGIT_SELECTION <= "01";
		SHIFT_SELECTION <= "000";
		WAIT FOR 20 ns;
		DIGIT_SELECTION <= "01";
		SHIFT_SELECTION <= "001";
		WAIT FOR 20 ns;
		DIGIT_SELECTION <= "10";
		SHIFT_SELECTION <= "011";
		WAIT FOR 20 ns;
		DIGIT_SELECTION <= "11";
		SHIFT_SELECTION <= "100";
		WAIT;
	END PROCESS;

	DUT : part2
	PORT MAP(SW(1 DOWNTO 0) => DIGIT_SELECTION,
		SW(4 DOWNTO 2) => SHIFT_SELECTION,
		HEX0 => DIG0,
		HEX1 => DIG1,
		HEX2 => DIG2,
		HEX3 => DIG3,
		HEX4 => DIG4);

END Behavior;